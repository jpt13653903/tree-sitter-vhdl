process(all) begin
  if    A1 then
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
  elsif A2 then
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
  elsif A3 then
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
  elsif A4 then
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
  elsif A5 then
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
  elsif A6 then
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
  elsif A7 then
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
  elsif A8 then
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
  elsif A9 then
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
  else
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
    A <= B;
  end if;
end process;

