================================================================================
Built-in libraries, operator overloading and a basic architecture body
================================================================================

library work;
    use work.whatnot.all;

library std;
    use std.whatnot.all;

library ieee;
    use ieee.whatnot.all;

entity Full_Adder is
  port(
    Clk   : in  std_logic;
    Reset : in  std_logic
  );
end entity Full_Adder;

-- A body of entity Full_Adder:
architecture DataFlow of Full_Adder is
  signal A, B: Bit;

  function "-"    (A : std_logic) return integer;
  function "??"   (A : std_logic) return integer;
  function "and"  (A : std_logic) return integer;
  function "or"   (A : std_logic) return integer;
  function "nand" (A : std_logic) return integer;
  function "nor"  (A : std_logic) return integer;
  function "xor"  (A : std_logic) return integer;
  function "xnor" (A : std_logic) return integer;
  function "="    (A : std_logic) return integer;
  function "/="   (A : std_logic) return integer;
  function "<"    (A : std_logic) return integer;
  function "<="   (A : std_logic) return integer;
  function ">"    (A : std_logic) return integer;
  function ">="   (A : std_logic) return integer;
  function "?="   (A : std_logic) return integer;
  function "?/="  (A : std_logic) return integer;
  function "?<"   (A : std_logic) return integer;
  function "?<="  (A : std_logic) return integer;
  function "?>"   (A : std_logic) return integer;
  function "?>="  (A : std_logic) return integer;
  function "sll"  (A : std_logic) return integer;
  function "srl"  (A : std_logic) return integer;
  function "sla"  (A : std_logic) return integer;
  function "sra"  (A : std_logic) return integer;
  function "rol"  (A : std_logic) return integer;
  function "ror"  (A : std_logic) return integer;
  function "+"    (A : std_logic) return integer;
  function "-"    (A : std_logic) return integer;
  function "&"    (A : std_logic) return integer;
  function "*"    (A : std_logic) return integer;
  function "/"    (A : std_logic) return integer;
  function "mod"  (A : std_logic) return integer;
  function "rem"  (A : std_logic) return integer;
  function "**"   (A : std_logic) return integer;
  function "abs"  (A : std_logic) return integer;
  function "not"  (A : std_logic) return integer;

  function MyFunc (A : std_logic) return integer;
begin
  MyInstance: entity work.Whatnot port map(
    Clock => Clk,
    Reset => Reset
  );

  A    <= X xor Y;
  B    <= A and Cin;
  Sum  <= A xor Cin;
  Cout <= B or (X and Y);

  process(A, B, C) is
    constant B : float := 8.291;
    variable A : integer := 5;
  begin
    if(rising_edge(Clk)) then
        A <= 5;
    else
        C <= 7;
    end if;
    for n in 0 to 3 loop
      case(WrRegisters.BenchTesting.HBW_Select(n)) is
        when "01"   => opHBW_SEL(n+1) <= '1';
        when "10"   => opHBW_SEL(n+1) <= '0';
        when others => opHBW_SEL(n+1) <= ipUSER_DIP(n);
      end case;
    end loop;
  end process;
  opHBW_SEL_N <= not(opHBW_SEL);
end architecture DataFlow;

--------------------------------------------------------------------------------

(design_file
  (design_unit
    (library_clause
      (LIBRARY)
      (logical_name_list
        (library_namespace))))
  (design_unit
    (use_clause
      (USE)
      (selected_name
        (library_namespace)
        (identifier)
        (ALL))))
  (design_unit
    (library_clause
      (LIBRARY)
      (logical_name_list
        (library_namespace))))
  (design_unit
    (use_clause
      (USE)
      (selected_name
        (library_namespace)
        (identifier)
        (ALL))))
  (design_unit
    (library_clause
      (LIBRARY)
      (logical_name_list
        (library_namespace))))
  (design_unit
    (use_clause
      (USE)
      (selected_name
        (library_namespace)
        (identifier)
        (ALL))))
  (design_unit
    (entity_declaration
      (ENTITY)
      (identifier)
      (entity_head
        (IS)
        (port_clause
          (PORT)
          (interface_list
            (interface_declaration
              (identifier_list
                (identifier))
              (simple_mode_indication
                (mode
                  (IN))
                (subtype_indication
                  (name
                    (library_type)))))
            (interface_declaration
              (identifier_list
                (identifier))
              (simple_mode_indication
                (mode
                  (IN))
                (subtype_indication
                  (name
                    (library_type))))))))
      (end_entity
        (END)
        (ENTITY)
        (identifier))))
  (comment)
  (design_unit
    (architecture_definition
      (ARCHITECTURE)
      (identifier)
      (OF)
      (name
        (identifier))
      (architecture_head
        (IS)
        (signal_declaration
          (SIGNAL)
          (identifier_list
            (identifier)
            (identifier))
          (subtype_indication
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (operator_symbol)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type))))
        (subprogram_declaration
          (function_specification
            (FUNCTION)
            (identifier)
            (parameter_list_specification
              (interface_list
                (interface_declaration
                  (identifier_list
                    (identifier))
                  (simple_mode_indication
                    (subtype_indication
                      (name
                        (library_type)))))))
            (RETURN)
            (name
              (library_type)))))
      (concurrent_block
        (BEGIN)
        (component_instantiation_statement
          (label_declaration
            (label))
          (instantiated_unit
            (ENTITY)
            (library_namespace)
            (name
              (identifier)))
          (port_map_aspect
            (PORT)
            (MAP)
            (association_list
              (association_element
                (name
                  (identifier))
                (conditional_expression
                  (simple_expression
                    (name
                      (identifier)))))
              (association_element
                (name
                  (identifier))
                (conditional_expression
                  (simple_expression
                    (name
                      (identifier))))))))
        (concurrent_simple_signal_assignment
          (name
            (identifier))
          (signal_assignment)
          (waveform
            (waveform_element
              (logical_expression
                (simple_expression
                  (name
                    (identifier)))
                (logical_operator)
                (simple_expression
                  (name
                    (identifier)))))))
        (concurrent_simple_signal_assignment
          (name
            (identifier))
          (signal_assignment)
          (waveform
            (waveform_element
              (logical_expression
                (simple_expression
                  (name
                    (identifier)))
                (logical_operator)
                (simple_expression
                  (name
                    (identifier)))))))
        (concurrent_simple_signal_assignment
          (name
            (identifier))
          (signal_assignment)
          (waveform
            (waveform_element
              (logical_expression
                (simple_expression
                  (name
                    (identifier)))
                (logical_operator)
                (simple_expression
                  (name
                    (identifier)))))))
        (concurrent_simple_signal_assignment
          (name
            (identifier))
          (signal_assignment)
          (waveform
            (waveform_element
              (logical_expression
                (simple_expression
                  (name
                    (identifier)))
                (logical_operator)
                (simple_expression
                  (parenthesis_expression
                    (element_association_list
                      (element_association
                        (conditional_expression
                          (logical_expression
                            (simple_expression
                              (name
                                (identifier)))
                            (logical_operator)
                            (simple_expression
                              (name
                                (identifier)))))))))))))
        (process_statement
          (PROCESS)
          (sensitivity_specification
            (sensitivity_list
              (name
                (identifier))
              (name
                (identifier))
              (name
                (identifier))))
          (process_head
            (IS)
            (constant_declaration
              (CONSTANT)
              (identifier_list
                (identifier))
              (subtype_indication
                (name
                  (library_type)))
              (initialiser
                (variable_assignment)
                (conditional_expression
                  (simple_expression
                    (decimal_literal_float)))))
            (variable_declaration
              (VARIABLE)
              (identifier_list
                (identifier))
              (subtype_indication
                (name
                  (library_type)))
              (initialiser
                (variable_assignment)
                (conditional_expression
                  (simple_expression
                    (decimal_literal))))))
          (sequential_block
            (BEGIN)
            (if_statement
              (if_expression
                (IF)
                (simple_expression
                  (parenthesis_expression
                    (element_association_list
                      (element_association
                        (conditional_expression
                          (simple_expression
                            (name
                              (library_function)
                              (name_selector
                                (parenthesis_group
                                  (association_or_range_list
                                    (association_element
                                      (conditional_expression
                                        (simple_expression
                                          (name
                                            (identifier))))))))))))))))
              (then_statements
                (THEN)
                (simple_waveform_assignment
                  (name
                    (identifier))
                  (signal_assignment)
                  (waveform
                    (waveform_element
                      (simple_expression
                        (decimal_literal))))))
              (else_statements
                (ELSE)
                (simple_waveform_assignment
                  (name
                    (identifier))
                  (signal_assignment)
                  (waveform
                    (waveform_element
                      (simple_expression
                        (decimal_literal))))))
              (end_if
                (END)
                (IF)))
            (loop_statement
              (for_loop
                (FOR)
                (parameter_specification
                  (identifier)
                  (IN)
                  (simple_range
                    (simple_expression
                      (decimal_literal))
                    (TO)
                    (simple_expression
                      (decimal_literal)))))
              (loop_body
                (LOOP)
                (case_statement
                  (case_expression
                    (CASE)
                    (simple_expression
                      (parenthesis_expression
                        (element_association_list
                          (element_association
                            (conditional_expression
                              (simple_expression
                                (name
                                  (identifier)
                                  (name_selector
                                    (selection
                                      (identifier)))
                                  (name_selector
                                    (selection
                                      (identifier)))
                                  (name_selector
                                    (parenthesis_group
                                      (association_or_range_list
                                        (association_element
                                          (conditional_expression
                                            (simple_expression
                                              (name
                                                (identifier))))))))))))))))
                  (case_body
                    (IS)
                    (case_statement_alternative
                      (when_element
                        (WHEN)
                        (simple_expression
                          (string_literal)))
                      (simple_waveform_assignment
                        (name
                          (identifier)
                          (name_selector
                            (parenthesis_group
                              (association_or_range_list
                                (association_element
                                  (conditional_expression
                                    (simple_expression
                                      (simple_expression
                                        (name
                                          (identifier)))
                                      (adding_operator)
                                      (simple_expression
                                        (decimal_literal)))))))))
                        (signal_assignment)
                        (waveform
                          (waveform_element
                            (simple_expression
                              (name
                                (library_constant_std_logic)))))))
                    (case_statement_alternative
                      (when_element
                        (WHEN)
                        (simple_expression
                          (string_literal)))
                      (simple_waveform_assignment
                        (name
                          (identifier)
                          (name_selector
                            (parenthesis_group
                              (association_or_range_list
                                (association_element
                                  (conditional_expression
                                    (simple_expression
                                      (simple_expression
                                        (name
                                          (identifier)))
                                      (adding_operator)
                                      (simple_expression
                                        (decimal_literal)))))))))
                        (signal_assignment)
                        (waveform
                          (waveform_element
                            (simple_expression
                              (name
                                (library_constant_std_logic)))))))
                    (case_statement_alternative
                      (when_element
                        (WHEN)
                        (OTHERS))
                      (simple_waveform_assignment
                        (name
                          (identifier)
                          (name_selector
                            (parenthesis_group
                              (association_or_range_list
                                (association_element
                                  (conditional_expression
                                    (simple_expression
                                      (simple_expression
                                        (name
                                          (identifier)))
                                      (adding_operator)
                                      (simple_expression
                                        (decimal_literal)))))))))
                        (signal_assignment)
                        (waveform
                          (waveform_element
                            (simple_expression
                              (name
                                (identifier)
                                (name_selector
                                  (parenthesis_group
                                    (association_or_range_list
                                      (association_element
                                        (conditional_expression
                                          (simple_expression
                                            (name
                                              (identifier)))))))))))))))
                  (end_case
                    (END)
                    (CASE))))
              (end_loop
                (END)
                (LOOP))))
          (end_process
            (END)
            (PROCESS)))
        (concurrent_simple_signal_assignment
          (name
            (identifier))
          (signal_assignment)
          (waveform
            (waveform_element
              (simple_expression
                (unary_operator)
                (simple_expression
                  (parenthesis_expression
                    (element_association_list
                      (element_association
                        (conditional_expression
                          (simple_expression
                            (name
                              (identifier)))))))))))))
      (end_architecture
        (END)
        (ARCHITECTURE)
        (identifier)))))

