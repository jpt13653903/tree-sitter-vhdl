MyLabel: if A1 generate
  A <= B;
elsif A2 generate
  A <= B;
elsif A3 generate
  A <= B;
elsif A4 generate
  A <= B;
elsif A5 generate
  A <= B;
elsif A6 generate
  A <= B;
elsif A7 generate
  A <= B;
elsif A8 generate
  A <= B;
elsif A9 generate
  A <= B;
else generate
  A <= B;
end generate;

